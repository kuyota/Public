module a();
  input wire a;
  input wire b;
  output wire c;


endmodule
